interface fa_intf;
  logic in1;
  logic in2;
  logic cin;
  logic sum, cout;
endinterface
